module ALUControl(
    wire input [1:0] ALUOp;
    wire input [5:0] functField;
    wire output [3:0] Operation;
)


always @(*) begin
    
end

